library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_unsigned.all;

package types is
  subtype opcodeT is std_logic_vector(5 downto 0);
  constant inop		: opcodeT := "000000";
  constant iadd		: opcodeT := "000001";
  constant isub		: opcodeT := "000100";
  constant ifneg	: opcodeT := "001111";
  constant iblt		: opcodeT := "010000";
  constant ibltf	: opcodeT := "010001";
  constant ibeq		: opcodeT := "010011";
  constant ibeqf	: opcodeT := "010100";
  constant ijmp		: opcodeT := "011110";
  constant ijmpr	: opcodeT := "100000";
  constant isave	: opcodeT := "100010";
  constant iseti1	: opcodeT := "100100";
  constant iseti2	: opcodeT := "100101";
  constant isetf1	: opcodeT := "100110";
  constant isetf2	: opcodeT := "100111";
  constant iload	: opcodeT := "101000";
  constant istore	: opcodeT := "101010";
  constant iinput	: opcodeT := "101100";
  constant iinputf	: opcodeT := "101101";
  constant ioutputint	: opcodeT := "110000";
  constant iloadb	: opcodeT := "110010";
  constant iloadbf	: opcodeT := "110011";
  constant istoreb	: opcodeT := "110100";
  constant istorebf	: opcodeT := "110101";
  constant iloadf	: opcodeT := "110110";
  constant istoref	: opcodeT := "110111";
  constant if2i		: opcodeT := "111001";
  constant iaddf	: opcodeT := "111010";
  constant isubf	: opcodeT := "111011";
  constant imulf	: opcodeT := "111100";
  constant iinvf	: opcodeT := "111101";
  constant isqrtf	: opcodeT := "111110";
  constant isli		: opcodeT := "111111";
end types;
